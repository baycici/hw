module ecc_encoder #(
	parameter DAT_WIDTH	=128,
	parameter ECC_WIDTH = 9
) (
    input   [DAT_WIDTH-1:0]   data_in, 
    output [ECC_WIDTH-1:0]   ecc_out
);

    wire [247:0] pattern [0:8];
	assign pattern[8] = 247'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	assign pattern[7] = 247'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
	assign pattern[6] = 247'b1111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111100000000000000000000000000;
	assign pattern[5] = 247'b1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000011111111111111100000000000;
	assign pattern[4] = 247'b1111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000111111110000000011111111000000001111111100000000111111110000000111111110000000011111111000000011111111000000011111110000;
	assign pattern[3] = 247'b1111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000111100001111000011110000111100001111000011110000111100001111000111100001111000011110000111100011110000111100011110001110;
	assign pattern[2] = 247'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110110011001100110011001100110011001100110011001100110011001100110110011001100110011001100110011011001100110011011001101101;
	assign pattern[1] = 247'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010110101010101010110101011011;
	assign pattern[0] = 247'b1001011001101001011010011001011001101001100101101001011001101001011010011001011010010110011010011001011001101001011010011001011011010011001011010010110011010011001011001101001011010011001011100101100110100101101001100101101101001100101110010110111;
    
    
    genvar i;
    generate
        for(i=0 ; i < ECC_WIDTH ; i=i+1)
            assign ecc_out[i] =   ^(data_in & pattern[i][DAT_WIDTH-1:0]);
    endgenerate
endmodule



