module ecc_decoder #(
	parameter DAT_WIDTH	=128,
	parameter ECC_WIDTH = 9
) (
    input   	[DAT_WIDTH-1:0]   	data_in, 
    input   	[ECC_WIDTH-1:0]   	ecc_in, 
	  output 	[DAT_WIDTH-1:0]		corrected_out,
    output  						single_error,
	  output						double_error,
	  output  						fault_error
);

  	reg [DAT_WIDTH-1:0] flip; 
    wire [ECC_WIDTH-1:0] check_bits, syndrome;  
    
    integer j, k;
    wire [247:0] pattern [0:8];
    // assign pattern[0] = 8'b11110000;
    // assign pattern[1] = 8'b10001110;
    // assign pattern[2] = 8'b01101101;
    // assign pattern[3] = 8'b01011011;
    // assign pattern[4] = 8'b10110111;
	assign pattern[8] = 247'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	assign pattern[7] = 247'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
	assign pattern[6] = 247'b1111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111100000000000000000000000000;
	assign pattern[5] = 247'b1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000011111111111111100000000000;
	assign pattern[4] = 247'b1111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000111111110000000011111111000000001111111100000000111111110000000111111110000000011111111000000011111111000000011111110000;
	assign pattern[3] = 247'b1111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000111100001111000011110000111100001111000011110000111100001111000111100001111000011110000111100011110000111100011110001110;
	assign pattern[2] = 247'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110110011001100110011001100110011001100110011001100110011001100110110011001100110011001100110011011001100110011011001101101;
	assign pattern[1] = 247'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010110101010101010110101011011;
	assign pattern[0] = 247'b1001011001101001011010011001011001101001100101101001011001101001011010011001011010010110011010011001011001101001011010011001011011010011001011010010110011010011001011001101001011010011001011100101100110100101101001100101101101001100101110010110111;

    genvar i;
    generate
        for(i=0 ; i < ECC_WIDTH ; i=i+1)
            assign check_bits[i] =   ^(data_in & pattern[i][DAT_WIDTH-1:0]);
    endgenerate

	assign syndrome = check_bits ^ ecc_in;
	
	always @(*)
	begin
		flip = {DAT_WIDTH{1'b1}};
		for(j=0;j<DAT_WIDTH;j=j+1)
		begin
			for(k=0;k<ECC_WIDTH;k=k+1)
			begin
				flip[j]= flip[j] & (~(syndrome[k]^pattern[k][j]));
			end
		end
	end
         
	assign corrected_out = flip ^ data_in;

	assign double_error = !(^syndrome) && |syndrome; //Even number of 1s in the signal syndrome, except for 0x0 
	assign single_error = |flip; 
	assign fault_error  = |(syndrome) && !double_error && !single_error ; 
	
endmodule
